module FanoutHash_37E9FE88073C5BAC (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  input logic [31:0] S7,
  input logic [31:0] S8,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
assign sel0 = (~E0) | (~S0[0]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[0]) | I2;
assign sel3 = (~E3) | (~S3[4]) | I3;
assign sel4 = (~E4) | (~S4[4]) | I4;
assign sel5 = (~E5) | (~S5[4]) | I5;
assign sel6 = (~E6) | (~S6[4]) | I6;
assign sel7 = (~E7) | (~S7[4]) | I7;
assign sel8 = (~E8) | (~S8[4]) | I8;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8;
endmodule   // FanoutHash_37E9FE88073C5BAC


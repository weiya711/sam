module FanoutHash_82899D6851EDC11 (
  input logic E0,
  input logic E1,
  input logic E10,
  input logic E11,
  input logic E12,
  input logic E13,
  input logic E14,
  input logic E15,
  input logic E16,
  input logic E17,
  input logic E18,
  input logic E19,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic E7,
  input logic E8,
  input logic E9,
  input logic I0,
  input logic I1,
  input logic I10,
  input logic I11,
  input logic I12,
  input logic I13,
  input logic I14,
  input logic I15,
  input logic I16,
  input logic I17,
  input logic I18,
  input logic I19,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic I7,
  input logic I8,
  input logic I9,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S10,
  input logic [7:0] S11,
  input logic [7:0] S12,
  input logic [7:0] S13,
  input logic [7:0] S14,
  input logic [7:0] S15,
  input logic [7:0] S16,
  input logic [7:0] S17,
  input logic [7:0] S18,
  input logic [7:0] S19,
  input logic [7:0] S2,
  input logic [7:0] S3,
  input logic [7:0] S4,
  input logic [7:0] S5,
  input logic [7:0] S6,
  input logic [7:0] S7,
  input logic [7:0] S8,
  input logic [7:0] S9,
  output logic O
);

logic sel0;
logic sel1;
logic sel10;
logic sel11;
logic sel12;
logic sel13;
logic sel14;
logic sel15;
logic sel16;
logic sel17;
logic sel18;
logic sel19;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
logic sel7;
logic sel8;
logic sel9;
assign sel0 = (~E0) | (~S0[4]) | I0;
assign sel1 = (~E1) | (~S1[4]) | I1;
assign sel2 = (~E2) | (~S2[4]) | I2;
assign sel3 = (~E3) | (~S3[4]) | I3;
assign sel4 = (~E4) | (~S4[4]) | I4;
assign sel5 = (~E5) | (~S5[4]) | I5;
assign sel6 = (~E6) | (~S6[4]) | I6;
assign sel7 = (~E7) | (~S7[4]) | I7;
assign sel8 = (~E8) | (~S8[4]) | I8;
assign sel9 = (~E9) | (~S9[4]) | I9;
assign sel10 = (~E10) | (~S10[4]) | I10;
assign sel11 = (~E11) | (~S11[4]) | I11;
assign sel12 = (~E12) | (~S12[4]) | I12;
assign sel13 = (~E13) | (~S13[4]) | I13;
assign sel14 = (~E14) | (~S14[4]) | I14;
assign sel15 = (~E15) | (~S15[4]) | I15;
assign sel16 = (~E16) | (~S16[4]) | I16;
assign sel17 = (~E17) | (~S17[4]) | I17;
assign sel18 = (~E18) | (~S18[4]) | I18;
assign sel19 = (~E19) | (~S19[4]) | I19;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6 & sel7 & sel8 & sel9 & sel10 &
    sel11 & sel12 & sel13 & sel14 & sel15 & sel16 & sel17 & sel18 & sel19;
endmodule   // FanoutHash_82899D6851EDC11


module FanoutHash_5D7AEC1255CDC1CC (
  input logic E0,
  input logic E1,
  input logic E2,
  input logic E3,
  input logic E4,
  input logic E5,
  input logic E6,
  input logic I0,
  input logic I1,
  input logic I2,
  input logic I3,
  input logic I4,
  input logic I5,
  input logic I6,
  input logic [7:0] S0,
  input logic [7:0] S1,
  input logic [7:0] S2,
  input logic [31:0] S3,
  input logic [31:0] S4,
  input logic [31:0] S5,
  input logic [31:0] S6,
  output logic O
);

logic sel0;
logic sel1;
logic sel2;
logic sel3;
logic sel4;
logic sel5;
logic sel6;
assign sel0 = (~E0) | (~S0[1]) | I0;
assign sel1 = (~E1) | (~S1[1]) | I1;
assign sel2 = (~E2) | (~S2[2]) | I2;
assign sel3 = (~E3) | (~S3[18]) | I3;
assign sel4 = (~E4) | (~S4[18]) | I4;
assign sel5 = (~E5) | (~S5[18]) | I5;
assign sel6 = (~E6) | (~S6[18]) | I6;
assign O = sel0 & sel1 & sel2 & sel3 & sel4 & sel5 & sel6;
endmodule   // FanoutHash_5D7AEC1255CDC1CC

